class axi4lite_test extends uvm_test;
  `uvm_component_utils(axi4lite_test)
  
  axi4lite_env env;
  
  function new(string name = "axi4lite_test", uvm_component parent);
    super.new(name, parent);
    `uvm_info("TEST_CLASS","Inside axi4lite_test constructor!", UVM_HIGH)
  endfunction: new
  
  function void build_phase(uvm_phase phase);
    super.build_phase(phase);
    `uvm_info("TEST_CLASS","Inside axi4lite_test build_phase!", UVM_HIGH)
    
    env = axi4lite_env::type_id::create("env",this);
    
  endfunction: build_phase
  
  function void connect_phase(uvm_phase phase);
     super.connect_phase(phase);
    `uvm_info("TEST_CLASS","Inside axi4lite_test connect_phase!", UVM_HIGH)
  endfunction: connect_phase
  
  task run_phase(uvm_phase phase);
    super.run_phase(phase);
    
    //Fill with logic later
    
  endtask: run_phase
  
endclass: axi4lite_test
